VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sutherland1989
  CLASS BLOCK ;
  FOREIGN sutherland1989 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.050 BY 0.050 ;
END sutherland1989
END LIBRARY

