VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NOR3
  CLASS CORE ;
  FOREIGN NOR3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.500 BY 5.050 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.800 4.500 5.300 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.250 4.500 0.250 ;
    END
  END VGND
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 0.350 0.850 0.750 0.900 ;
        RECT 2.600 0.850 3.000 0.900 ;
        RECT 0.350 0.550 3.000 0.850 ;
        RECT 0.350 0.500 0.750 0.550 ;
        RECT 2.600 0.500 3.000 0.550 ;
    END
  END Y
  PIN A1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 2.050 2.400 2.450 3.200 ;
    END
  END A1
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 0.950 2.400 1.300 3.200 ;
    END
  END A
  PIN A2
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 3.150 2.400 3.550 3.200 ;
    END
  END A2
END NOR3
END LIBRARY

