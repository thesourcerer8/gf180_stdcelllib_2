MACRO AAAOAI3322
 CLASS CORE ;
 FOREIGN AAAOAI3322 0 0 ;
 SIZE 13.44 BY 5.04 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 4.80000000 13.44000000 5.28000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 13.44000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.37000000 3.20700000 0.75000000 3.25700000 ;
        RECT 2.61000000 3.20700000 2.99000000 3.25700000 ;
        RECT 0.37000000 3.25700000 2.99000000 3.53700000 ;
        RECT 0.37000000 3.53700000 0.75000000 3.58700000 ;
        RECT 2.61000000 3.53700000 2.99000000 3.58700000 ;
    END
  END Y

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 4.29000000 2.39700000 4.67000000 2.77700000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 5.41000000 2.39700000 5.79000000 2.77700000 ;
    END
  END B1

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 2.05000000 2.39700000 2.43000000 2.77700000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 3.17000000 2.39700000 3.55000000 2.77700000 ;
    END
  END A2

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 6.53000000 2.39700000 6.91000000 2.77700000 ;
    END
  END B

  PIN D1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 9.89000000 2.80200000 10.27000000 3.18200000 ;
    END
  END D1

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 8.77000000 2.80200000 9.15000000 3.18200000 ;
    END
  END D

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 11.01000000 3.07200000 11.39000000 3.45200000 ;
    END
  END C1

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 7.70000000 2.17700000 11.90000000 2.39700000 ;
        RECT 7.70000000 2.39700000 11.95000000 2.45700000 ;
        RECT 11.57000000 2.45700000 11.95000000 2.77700000 ;
        RECT 7.70000000 2.45700000 7.98000000 2.80200000 ;
        RECT 7.65000000 2.80200000 8.03000000 3.18200000 ;
    END
  END C

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.93000000 2.39700000 1.31000000 2.77700000 ;
    END
  END A

 OBS
    LAYER polycont ;
     RECT 1.01000000 2.47700000 1.23000000 2.69700000 ;
     RECT 2.13000000 2.47700000 2.35000000 2.69700000 ;
     RECT 3.25000000 2.47700000 3.47000000 2.69700000 ;
     RECT 4.37000000 2.47700000 4.59000000 2.69700000 ;
     RECT 5.49000000 2.47700000 5.71000000 2.69700000 ;
     RECT 6.61000000 2.47700000 6.83000000 2.69700000 ;
     RECT 8.85000000 2.47700000 9.07000000 2.69700000 ;
     RECT 9.97000000 2.47700000 10.19000000 2.69700000 ;
     RECT 11.09000000 2.47700000 11.31000000 2.69700000 ;
     RECT 12.21000000 2.47700000 12.43000000 2.69700000 ;
     RECT 1.01000000 2.88200000 1.23000000 3.10200000 ;
     RECT 2.13000000 2.88200000 2.35000000 3.10200000 ;
     RECT 3.25000000 2.88200000 3.47000000 3.10200000 ;
     RECT 4.37000000 2.88200000 4.59000000 3.10200000 ;
     RECT 5.49000000 2.88200000 5.71000000 3.10200000 ;
     RECT 6.61000000 2.88200000 6.83000000 3.10200000 ;
     RECT 7.73000000 2.88200000 7.95000000 3.10200000 ;
     RECT 8.85000000 2.88200000 9.07000000 3.10200000 ;
     RECT 9.97000000 2.88200000 10.19000000 3.10200000 ;
     RECT 11.09000000 2.88200000 11.31000000 3.10200000 ;

    LAYER pdiffc ;
     RECT 0.45000000 3.28700000 0.67000000 3.50700000 ;
     RECT 2.69000000 3.28700000 2.91000000 3.50700000 ;
     RECT 3.81000000 3.28700000 4.03000000 3.50700000 ;
     RECT 6.05000000 3.28700000 6.27000000 3.50700000 ;
     RECT 8.29000000 3.28700000 8.51000000 3.64200000 ;
     RECT 10.53000000 3.42200000 10.75000000 3.64200000 ;
     RECT 4.93000000 3.82700000 5.15000000 4.04700000 ;
     RECT 7.17000000 3.82700000 7.39000000 4.04700000 ;
     RECT 11.65000000 3.82700000 11.87000000 4.04700000 ;
     RECT 1.57000000 4.09700000 1.79000000 4.31700000 ;
     RECT 9.41000000 4.50200000 9.63000000 4.72200000 ;

    LAYER ndiffc ;
     RECT 3.81000000 0.31700000 4.03000000 0.53700000 ;
     RECT 10.53000000 0.31700000 10.75000000 0.53700000 ;
     RECT 7.17000000 1.39700000 7.39000000 1.61700000 ;
     RECT 0.45000000 1.93700000 0.67000000 2.15700000 ;
     RECT 8.29000000 1.93700000 8.51000000 2.15700000 ;
     RECT 12.77000000 1.93700000 12.99000000 2.15700000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 13.44000000 0.24000000 ;
     RECT 3.73000000 0.24000000 4.11000000 0.61700000 ;
     RECT 10.45000000 0.24000000 10.83000000 0.61700000 ;
     RECT 7.09000000 1.31700000 7.47000000 1.69700000 ;
     RECT 12.69000000 1.85700000 13.07000000 2.23700000 ;
     RECT 11.57000000 2.39700000 11.95000000 2.47200000 ;
     RECT 12.13000000 2.39700000 12.51000000 2.47200000 ;
     RECT 11.57000000 2.47200000 12.51000000 2.70200000 ;
     RECT 11.57000000 2.70200000 11.95000000 2.77700000 ;
     RECT 12.13000000 2.70200000 12.51000000 2.77700000 ;
     RECT 0.93000000 2.39700000 1.31000000 3.18200000 ;
     RECT 2.05000000 2.39700000 2.43000000 3.18200000 ;
     RECT 3.17000000 2.39700000 3.55000000 3.18200000 ;
     RECT 4.29000000 2.39700000 4.67000000 3.18200000 ;
     RECT 5.41000000 2.39700000 5.79000000 3.18200000 ;
     RECT 6.53000000 2.39700000 6.91000000 3.18200000 ;
     RECT 7.65000000 2.80200000 8.03000000 3.18200000 ;
     RECT 8.77000000 2.39700000 9.15000000 3.18200000 ;
     RECT 9.89000000 2.39700000 10.27000000 3.18200000 ;
     RECT 11.01000000 2.39700000 11.39000000 3.45200000 ;
     RECT 0.37000000 1.85700000 0.75000000 2.23700000 ;
     RECT 0.44500000 2.23700000 0.67500000 3.20700000 ;
     RECT 0.37000000 3.20700000 0.75000000 3.58700000 ;
     RECT 2.61000000 3.20700000 2.99000000 3.58700000 ;
     RECT 3.73000000 3.20700000 4.11000000 3.58700000 ;
     RECT 5.97000000 1.31700000 6.35000000 1.69700000 ;
     RECT 6.04500000 1.69700000 6.27500000 3.07200000 ;
     RECT 5.97000000 3.07200000 6.35000000 3.58700000 ;
     RECT 8.21000000 1.85700000 8.59000000 2.23700000 ;
     RECT 8.28500000 2.23700000 8.51500000 3.20700000 ;
     RECT 8.21000000 3.20700000 8.59000000 3.41700000 ;
     RECT 10.45000000 3.34200000 10.83000000 3.41700000 ;
     RECT 8.21000000 3.41700000 10.83000000 3.64700000 ;
     RECT 8.21000000 3.64700000 8.59000000 3.72200000 ;
     RECT 10.45000000 3.64700000 10.83000000 3.72200000 ;
     RECT 4.85000000 3.74700000 5.23000000 4.12700000 ;
     RECT 7.09000000 3.74700000 7.47000000 4.12700000 ;
     RECT 11.57000000 3.74700000 11.95000000 4.12700000 ;
     RECT 1.49000000 4.01700000 1.87000000 4.39700000 ;
     RECT 9.33000000 4.42200000 9.71000000 4.80000000 ;
     RECT 0.00000000 4.80000000 13.44000000 5.28000000 ;

    LAYER via1 ;
     RECT 6.03000000 1.37700000 6.29000000 1.63700000 ;
     RECT 7.15000000 1.37700000 7.41000000 1.63700000 ;
     RECT 12.75000000 1.91700000 13.01000000 2.17700000 ;
     RECT 0.99000000 2.45700000 1.25000000 2.71700000 ;
     RECT 2.11000000 2.45700000 2.37000000 2.71700000 ;
     RECT 3.23000000 2.45700000 3.49000000 2.71700000 ;
     RECT 4.35000000 2.45700000 4.61000000 2.71700000 ;
     RECT 5.47000000 2.45700000 5.73000000 2.71700000 ;
     RECT 6.59000000 2.45700000 6.85000000 2.71700000 ;
     RECT 11.63000000 2.45700000 11.89000000 2.71700000 ;
     RECT 7.71000000 2.86200000 7.97000000 3.12200000 ;
     RECT 8.83000000 2.86200000 9.09000000 3.12200000 ;
     RECT 9.95000000 2.86200000 10.21000000 3.12200000 ;
     RECT 6.03000000 3.13200000 6.29000000 3.39200000 ;
     RECT 11.07000000 3.13200000 11.33000000 3.39200000 ;
     RECT 0.43000000 3.26700000 0.69000000 3.52700000 ;
     RECT 2.67000000 3.26700000 2.93000000 3.52700000 ;
     RECT 3.79000000 3.26700000 4.05000000 3.52700000 ;
     RECT 4.91000000 3.80700000 5.17000000 4.06700000 ;
     RECT 7.15000000 3.80700000 7.41000000 4.06700000 ;
     RECT 11.63000000 3.80700000 11.89000000 4.06700000 ;
     RECT 1.55000000 4.07700000 1.81000000 4.33700000 ;

    LAYER met2 ;
     RECT 5.97000000 1.31700000 6.35000000 1.36700000 ;
     RECT 7.09000000 1.31700000 7.47000000 1.36700000 ;
     RECT 5.97000000 1.36700000 7.47000000 1.64700000 ;
     RECT 5.97000000 1.64700000 6.35000000 1.69700000 ;
     RECT 7.09000000 1.64700000 7.47000000 1.69700000 ;
     RECT 0.93000000 2.39700000 1.31000000 2.77700000 ;
     RECT 2.05000000 2.39700000 2.43000000 2.77700000 ;
     RECT 3.17000000 2.39700000 3.55000000 2.77700000 ;
     RECT 4.29000000 2.39700000 4.67000000 2.77700000 ;
     RECT 5.41000000 2.39700000 5.79000000 2.77700000 ;
     RECT 6.53000000 2.39700000 6.91000000 2.77700000 ;
     RECT 7.70000000 2.17700000 11.90000000 2.39700000 ;
     RECT 7.70000000 2.39700000 11.95000000 2.45700000 ;
     RECT 11.57000000 2.45700000 11.95000000 2.77700000 ;
     RECT 7.70000000 2.45700000 7.98000000 2.80200000 ;
     RECT 7.65000000 2.80200000 8.03000000 3.18200000 ;
     RECT 8.77000000 2.80200000 9.15000000 3.18200000 ;
     RECT 9.89000000 2.80200000 10.27000000 3.18200000 ;
     RECT 11.01000000 3.07200000 11.39000000 3.45200000 ;
     RECT 0.37000000 3.20700000 0.75000000 3.25700000 ;
     RECT 2.61000000 3.20700000 2.99000000 3.25700000 ;
     RECT 0.37000000 3.25700000 2.99000000 3.53700000 ;
     RECT 0.37000000 3.53700000 0.75000000 3.58700000 ;
     RECT 2.61000000 3.53700000 2.99000000 3.58700000 ;
     RECT 12.69000000 1.85700000 13.07000000 2.23700000 ;
     RECT 4.85000000 3.74700000 5.23000000 3.79700000 ;
     RECT 7.09000000 3.74700000 7.47000000 3.79700000 ;
     RECT 11.57000000 3.74700000 11.95000000 3.79700000 ;
     RECT 12.74000000 2.23700000 13.02000000 3.79700000 ;
     RECT 4.85000000 3.79700000 13.02000000 4.07700000 ;
     RECT 4.85000000 4.07700000 5.23000000 4.12700000 ;
     RECT 7.09000000 4.07700000 7.47000000 4.12700000 ;
     RECT 11.57000000 4.07700000 11.95000000 4.12700000 ;
     RECT 5.97000000 3.07200000 6.35000000 3.12200000 ;
     RECT 3.78000000 3.12200000 6.35000000 3.20700000 ;
     RECT 3.73000000 3.20700000 6.35000000 3.40200000 ;
     RECT 5.97000000 3.40200000 6.35000000 3.45200000 ;
     RECT 3.73000000 3.40200000 4.11000000 3.58700000 ;
     RECT 1.49000000 4.01700000 1.87000000 4.06700000 ;
     RECT 3.78000000 3.58700000 4.06000000 4.06700000 ;
     RECT 1.49000000 4.06700000 4.06000000 4.34700000 ;
     RECT 1.49000000 4.34700000 1.87000000 4.39700000 ;

 END
END AAAOAI3322
