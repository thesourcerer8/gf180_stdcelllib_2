MACRO VANBERKEL1991
 CLASS CORE ;
 FOREIGN VANBERKEL1991 0 0 ;
 SIZE 8.96 BY 5.04 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 4.80000000 8.96000000 5.28000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 8.96000000 0.24000000 ;
    END
  END GND

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 5.41000000 1.58700000 5.79000000 1.63700000 ;
        RECT 8.21000000 1.58700000 8.59000000 1.63700000 ;
        RECT 5.41000000 1.63700000 8.59000000 1.91700000 ;
        RECT 5.41000000 1.91700000 5.79000000 1.96700000 ;
        RECT 8.21000000 1.91700000 8.59000000 1.96700000 ;
    END
  END C

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 3.17000000 1.58700000 3.55000000 1.63700000 ;
        RECT 0.98000000 1.63700000 3.55000000 1.91700000 ;
        RECT 3.17000000 1.91700000 3.55000000 1.96700000 ;
        RECT 0.98000000 1.91700000 1.26000000 2.39700000 ;
        RECT 0.93000000 2.39700000 1.31000000 3.18200000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 2.05000000 2.39700000 2.43000000 2.85200000 ;
        RECT 6.53000000 2.39700000 6.91000000 2.85200000 ;
        RECT 2.05000000 2.85200000 6.91000000 3.13200000 ;
        RECT 2.05000000 3.13200000 2.43000000 3.18200000 ;
        RECT 6.53000000 3.13200000 6.91000000 3.18200000 ;
    END
  END A

 OBS
    LAYER polycont ;
     RECT 1.01000000 2.47700000 1.23000000 2.69700000 ;
     RECT 2.13000000 2.47700000 2.35000000 2.69700000 ;
     RECT 3.25000000 2.47700000 3.47000000 2.69700000 ;
     RECT 5.49000000 2.47700000 5.71000000 2.69700000 ;
     RECT 6.61000000 2.47700000 6.83000000 2.69700000 ;
     RECT 7.73000000 2.47700000 7.95000000 2.69700000 ;
     RECT 1.01000000 2.88200000 1.23000000 3.10200000 ;
     RECT 2.13000000 2.88200000 2.35000000 3.10200000 ;
     RECT 3.25000000 2.88200000 3.47000000 3.10200000 ;
     RECT 5.49000000 2.88200000 5.71000000 3.10200000 ;
     RECT 6.61000000 2.88200000 6.83000000 3.10200000 ;
     RECT 7.73000000 2.88200000 7.95000000 3.10200000 ;

    LAYER pdiffc ;
     RECT 1.57000000 3.28700000 1.79000000 3.50700000 ;
     RECT 8.29000000 3.28700000 8.51000000 3.50700000 ;
     RECT 2.69000000 3.42200000 2.91000000 3.64200000 ;
     RECT 4.93000000 3.42200000 5.15000000 3.64200000 ;
     RECT 1.57000000 3.55700000 1.79000000 3.77700000 ;
     RECT 0.45000000 4.23200000 0.67000000 4.45200000 ;
     RECT 6.05000000 4.23200000 6.27000000 4.45200000 ;
     RECT 3.81000000 4.50200000 4.03000000 4.72200000 ;
     RECT 7.17000000 4.50200000 7.39000000 4.72200000 ;

    LAYER ndiffc ;
     RECT 3.81000000 0.31700000 4.03000000 0.53700000 ;
     RECT 7.17000000 0.31700000 7.39000000 0.53700000 ;
     RECT 0.45000000 0.58700000 0.67000000 0.80700000 ;
     RECT 6.05000000 0.58700000 6.27000000 0.80700000 ;
     RECT 2.69000000 0.85700000 2.91000000 1.07700000 ;
     RECT 4.93000000 0.85700000 5.15000000 1.07700000 ;
     RECT 8.29000000 1.66700000 8.51000000 1.88700000 ;
     RECT 1.57000000 1.93700000 1.79000000 2.15700000 ;
     RECT 8.29000000 1.93700000 8.51000000 2.15700000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 8.96000000 0.24000000 ;
     RECT 3.73000000 0.24000000 4.11000000 0.61700000 ;
     RECT 7.09000000 0.24000000 7.47000000 0.61700000 ;
     RECT 0.37000000 0.50700000 0.75000000 0.88700000 ;
     RECT 5.97000000 0.50700000 6.35000000 0.88700000 ;
     RECT 2.61000000 0.77700000 2.99000000 0.85200000 ;
     RECT 4.85000000 0.77700000 5.23000000 0.85200000 ;
     RECT 2.61000000 0.85200000 5.23000000 1.08200000 ;
     RECT 2.61000000 1.08200000 2.99000000 1.15700000 ;
     RECT 4.85000000 1.08200000 5.23000000 1.15700000 ;
     RECT 0.93000000 2.39700000 1.31000000 2.77700000 ;
     RECT 2.05000000 2.39700000 2.43000000 2.77700000 ;
     RECT 6.53000000 2.39700000 6.91000000 2.77700000 ;
     RECT 7.65000000 2.39700000 8.03000000 2.77700000 ;
     RECT 0.93000000 2.80200000 1.31000000 3.18200000 ;
     RECT 2.05000000 2.80200000 2.43000000 3.18200000 ;
     RECT 3.17000000 1.58700000 3.55000000 1.96700000 ;
     RECT 3.24500000 1.96700000 3.47500000 2.39700000 ;
     RECT 3.17000000 2.39700000 3.55000000 3.18200000 ;
     RECT 5.41000000 1.58700000 5.79000000 1.96700000 ;
     RECT 5.48500000 1.96700000 5.71500000 2.39700000 ;
     RECT 5.41000000 2.39700000 5.79000000 3.18200000 ;
     RECT 6.53000000 2.80200000 6.91000000 3.18200000 ;
     RECT 7.65000000 2.80200000 8.03000000 3.18200000 ;
     RECT 8.21000000 1.58700000 8.59000000 2.23700000 ;
     RECT 8.28500000 2.23700000 8.51500000 3.20700000 ;
     RECT 8.21000000 3.20700000 8.59000000 3.58700000 ;
     RECT 2.61000000 3.34200000 2.99000000 3.41700000 ;
     RECT 4.85000000 3.34200000 5.23000000 3.41700000 ;
     RECT 2.61000000 3.41700000 5.23000000 3.64700000 ;
     RECT 2.61000000 3.64700000 2.99000000 3.72200000 ;
     RECT 4.85000000 3.64700000 5.23000000 3.72200000 ;
     RECT 1.49000000 1.85700000 1.87000000 2.23700000 ;
     RECT 1.56500000 2.23700000 1.79500000 3.20700000 ;
     RECT 1.49000000 3.20700000 1.87000000 3.85700000 ;
     RECT 0.37000000 4.15200000 0.75000000 4.53200000 ;
     RECT 5.97000000 4.15200000 6.35000000 4.53200000 ;
     RECT 3.73000000 4.42200000 4.11000000 4.80000000 ;
     RECT 7.09000000 4.42200000 7.47000000 4.80000000 ;
     RECT 0.00000000 4.80000000 8.96000000 5.28000000 ;

    LAYER via1 ;
     RECT 0.43000000 0.56700000 0.69000000 0.82700000 ;
     RECT 6.03000000 0.56700000 6.29000000 0.82700000 ;
     RECT 3.23000000 1.64700000 3.49000000 1.90700000 ;
     RECT 5.47000000 1.64700000 5.73000000 1.90700000 ;
     RECT 8.27000000 1.64700000 8.53000000 1.90700000 ;
     RECT 0.99000000 2.45700000 1.25000000 2.71700000 ;
     RECT 2.11000000 2.45700000 2.37000000 2.71700000 ;
     RECT 6.59000000 2.45700000 6.85000000 2.71700000 ;
     RECT 7.71000000 2.45700000 7.97000000 2.71700000 ;
     RECT 0.99000000 2.86200000 1.25000000 3.12200000 ;
     RECT 2.11000000 2.86200000 2.37000000 3.12200000 ;
     RECT 6.59000000 2.86200000 6.85000000 3.12200000 ;
     RECT 7.71000000 2.86200000 7.97000000 3.12200000 ;
     RECT 1.55000000 3.53700000 1.81000000 3.79700000 ;
     RECT 0.43000000 4.21200000 0.69000000 4.47200000 ;
     RECT 6.03000000 4.21200000 6.29000000 4.47200000 ;

    LAYER met2 ;
     RECT 0.37000000 0.50700000 0.75000000 0.55700000 ;
     RECT 5.97000000 0.50700000 6.35000000 0.55700000 ;
     RECT 0.37000000 0.55700000 6.35000000 0.83700000 ;
     RECT 0.37000000 0.83700000 0.75000000 0.88700000 ;
     RECT 5.97000000 0.83700000 6.35000000 0.88700000 ;
     RECT 5.41000000 1.58700000 5.79000000 1.63700000 ;
     RECT 8.21000000 1.58700000 8.59000000 1.63700000 ;
     RECT 5.41000000 1.63700000 8.59000000 1.91700000 ;
     RECT 5.41000000 1.91700000 5.79000000 1.96700000 ;
     RECT 8.21000000 1.91700000 8.59000000 1.96700000 ;
     RECT 3.17000000 1.58700000 3.55000000 1.63700000 ;
     RECT 0.98000000 1.63700000 3.55000000 1.91700000 ;
     RECT 3.17000000 1.91700000 3.55000000 1.96700000 ;
     RECT 0.98000000 1.91700000 1.26000000 2.39700000 ;
     RECT 0.93000000 2.39700000 1.31000000 3.18200000 ;
     RECT 2.05000000 2.39700000 2.43000000 2.85200000 ;
     RECT 6.53000000 2.39700000 6.91000000 2.85200000 ;
     RECT 2.05000000 2.85200000 6.91000000 3.13200000 ;
     RECT 2.05000000 3.13200000 2.43000000 3.18200000 ;
     RECT 6.53000000 3.13200000 6.91000000 3.18200000 ;
     RECT 7.65000000 2.39700000 8.03000000 3.18200000 ;
     RECT 1.49000000 3.47700000 1.87000000 3.52700000 ;
     RECT 7.70000000 3.18200000 7.98000000 3.52700000 ;
     RECT 1.49000000 3.52700000 7.98000000 3.80700000 ;
     RECT 1.49000000 3.80700000 1.87000000 3.85700000 ;
     RECT 0.37000000 4.15200000 0.75000000 4.20200000 ;
     RECT 5.97000000 4.15200000 6.35000000 4.20200000 ;
     RECT 0.37000000 4.20200000 6.35000000 4.48200000 ;
     RECT 0.37000000 4.48200000 0.75000000 4.53200000 ;
     RECT 5.97000000 4.48200000 6.35000000 4.53200000 ;

 END
END VANBERKEL1991
