MACRO NOR3
 CLASS CORE ;
 FOREIGN NOR3 0 0 ;
 SIZE 4.48 BY 5.04 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 4.80000000 4.48000000 5.28000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 4.48000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.37000000 0.50700000 0.75000000 0.55700000 ;
        RECT 2.61000000 0.50700000 2.99000000 0.55700000 ;
        RECT 0.37000000 0.55700000 2.99000000 0.83700000 ;
        RECT 0.37000000 0.83700000 0.75000000 0.88700000 ;
        RECT 2.61000000 0.83700000 2.99000000 0.88700000 ;
    END
  END Y

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 2.05000000 2.39700000 2.43000000 3.18200000 ;
    END
  END A1

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.93000000 2.39700000 1.31000000 3.18200000 ;
    END
  END A

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 3.17000000 2.39700000 3.55000000 3.18200000 ;
    END
  END A2

 OBS
    LAYER polycont ;
     RECT 1.01000000 2.47700000 1.23000000 2.69700000 ;
     RECT 2.13000000 2.47700000 2.35000000 2.69700000 ;
     RECT 3.25000000 2.47700000 3.47000000 2.69700000 ;
     RECT 1.01000000 2.88200000 1.23000000 3.10200000 ;
     RECT 2.13000000 2.88200000 2.35000000 3.10200000 ;
     RECT 3.25000000 2.88200000 3.47000000 3.10200000 ;

    LAYER pdiffc ;
     RECT 0.45000000 3.28700000 0.67000000 3.50700000 ;
     RECT 3.81000000 4.50200000 4.03000000 4.72200000 ;

    LAYER ndiffc ;
     RECT 1.57000000 0.31700000 1.79000000 0.53700000 ;
     RECT 3.81000000 0.31700000 4.03000000 0.53700000 ;
     RECT 0.45000000 0.58700000 0.67000000 0.80700000 ;
     RECT 2.69000000 0.58700000 2.91000000 0.80700000 ;
     RECT 0.45000000 1.93700000 0.67000000 2.15700000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 4.48000000 0.24000000 ;
     RECT 1.49000000 0.24000000 1.87000000 0.61700000 ;
     RECT 3.73000000 0.24000000 4.11000000 0.61700000 ;
     RECT 0.37000000 0.50700000 0.75000000 0.88700000 ;
     RECT 2.61000000 0.50700000 2.99000000 0.88700000 ;
     RECT 0.93000000 2.39700000 1.31000000 2.77700000 ;
     RECT 2.05000000 2.39700000 2.43000000 2.77700000 ;
     RECT 3.17000000 2.39700000 3.55000000 2.77700000 ;
     RECT 0.93000000 2.80200000 1.31000000 3.18200000 ;
     RECT 2.05000000 2.80200000 2.43000000 3.18200000 ;
     RECT 3.17000000 2.80200000 3.55000000 3.18200000 ;
     RECT 0.37000000 1.85700000 0.75000000 2.23700000 ;
     RECT 0.44500000 2.23700000 0.67500000 3.20700000 ;
     RECT 0.37000000 3.20700000 0.75000000 3.58700000 ;
     RECT 3.73000000 4.42200000 4.11000000 4.80000000 ;
     RECT 0.00000000 4.80000000 4.48000000 5.28000000 ;

    LAYER via1 ;
     RECT 0.43000000 0.56700000 0.69000000 0.82700000 ;
     RECT 2.67000000 0.56700000 2.93000000 0.82700000 ;
     RECT 0.99000000 2.45700000 1.25000000 2.71700000 ;
     RECT 2.11000000 2.45700000 2.37000000 2.71700000 ;
     RECT 3.23000000 2.45700000 3.49000000 2.71700000 ;
     RECT 0.99000000 2.86200000 1.25000000 3.12200000 ;
     RECT 2.11000000 2.86200000 2.37000000 3.12200000 ;
     RECT 3.23000000 2.86200000 3.49000000 3.12200000 ;

    LAYER met2 ;
     RECT 0.37000000 0.50700000 0.75000000 0.55700000 ;
     RECT 2.61000000 0.50700000 2.99000000 0.55700000 ;
     RECT 0.37000000 0.55700000 2.99000000 0.83700000 ;
     RECT 0.37000000 0.83700000 0.75000000 0.88700000 ;
     RECT 2.61000000 0.83700000 2.99000000 0.88700000 ;
     RECT 0.93000000 2.39700000 1.31000000 3.18200000 ;
     RECT 2.05000000 2.39700000 2.43000000 3.18200000 ;
     RECT 3.17000000 2.39700000 3.55000000 3.18200000 ;

 END
END NOR3
