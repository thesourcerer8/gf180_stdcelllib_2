VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vanberkel1991
  CLASS BLOCK ;
  FOREIGN vanberkel1991 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.050 BY 0.050 ;
END vanberkel1991
END LIBRARY

