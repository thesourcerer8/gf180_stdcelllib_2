VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OAAOAOI21311
  CLASS CORE ;
  FOREIGN OAAOAOI21311 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.300 BY 5.050 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.800 12.300 5.300 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.250 12.300 0.250 ;
    END
  END VGND
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 0.350 2.050 0.750 2.100 ;
        RECT 1.500 2.050 1.850 2.100 ;
        RECT 0.350 1.750 1.850 2.050 ;
        RECT 0.350 1.700 0.750 1.750 ;
        RECT 1.500 1.700 1.850 1.750 ;
    END
  END Y
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 4.300 2.400 4.650 2.800 ;
    END
  END B
  PIN C1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 6.550 2.400 6.900 2.800 ;
    END
  END C1
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 8.750 2.750 9.150 2.800 ;
        RECT 9.900 2.750 10.250 3.050 ;
        RECT 8.750 2.650 10.250 2.750 ;
        RECT 8.750 2.450 10.200 2.650 ;
        RECT 8.750 2.400 9.150 2.450 ;
    END
  END D
  PIN E
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 11.000 2.400 11.400 2.800 ;
    END
  END E
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 0.950 2.400 1.300 3.200 ;
    END
  END A
  PIN C2
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 7.650 2.400 8.050 2.800 ;
    END
  END C2
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 5.400 2.400 5.800 2.800 ;
    END
  END C
  PIN A1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 2.050 2.800 2.450 3.200 ;
    END
  END A1
END OAAOAOI21311
END LIBRARY

