VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO AAAOAOI33211
  CLASS CORE ;
  FOREIGN AAAOAOI33211 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.450 BY 5.050 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.800 13.450 5.300 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.250 13.450 0.250 ;
    END
  END VGND
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 0.350 3.400 0.750 3.450 ;
        RECT 2.600 3.400 3.000 3.450 ;
        RECT 0.350 3.100 3.000 3.400 ;
        RECT 0.350 3.050 0.750 3.100 ;
        RECT 2.600 3.050 3.000 3.100 ;
    END
  END Y
  PIN A2
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 3.150 2.400 3.550 2.800 ;
    END
  END A2
  PIN C1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 7.650 2.450 8.050 2.500 ;
        RECT 9.900 2.450 10.250 2.800 ;
        RECT 7.650 2.400 10.250 2.450 ;
        RECT 7.650 2.200 10.200 2.400 ;
        RECT 7.650 2.150 8.050 2.200 ;
    END
  END C1
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 0.950 2.400 1.300 2.800 ;
    END
  END A
  PIN B2
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 4.300 2.400 4.650 2.800 ;
    END
  END B2
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 8.750 2.800 9.150 3.200 ;
    END
  END C
  PIN E
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 12.150 2.400 12.500 2.800 ;
    END
  END E
  PIN B1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 5.400 2.400 5.800 2.800 ;
    END
  END B1
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 11.000 2.400 11.400 2.800 ;
    END
  END D
  PIN A1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 2.050 2.400 2.450 2.800 ;
    END
  END A1
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 6.550 2.400 6.900 2.800 ;
    END
  END B
END AAAOAOI33211
END LIBRARY

