MACRO OAI41
 CLASS CORE ;
 FOREIGN OAI41 0 0 ;
 SIZE 6.72 BY 5.04 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 4.80000000 6.72000000 5.28000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 6.72000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 2.61000000 0.50700000 2.99000000 0.55700000 ;
        RECT 4.85000000 0.50700000 5.23000000 0.55700000 ;
        RECT 2.61000000 0.55700000 5.23000000 0.83700000 ;
        RECT 2.61000000 0.83700000 2.99000000 0.88700000 ;
        RECT 4.85000000 0.83700000 5.23000000 0.88700000 ;
    END
  END Y

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 4.29000000 2.80200000 4.67000000 3.18200000 ;
    END
  END A1

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 1.49000000 2.39700000 1.87000000 2.77700000 ;
    END
  END B

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 1.49000000 3.07200000 1.87000000 3.45200000 ;
    END
  END A3

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 5.41000000 2.39700000 5.79000000 3.18200000 ;
    END
  END A

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 3.73000000 2.12700000 4.11000000 2.50700000 ;
    END
  END A2

 OBS
    LAYER polycont ;
     RECT 1.01000000 2.47700000 1.23000000 2.69700000 ;
     RECT 2.13000000 2.47700000 2.35000000 2.69700000 ;
     RECT 3.25000000 2.47700000 3.47000000 2.69700000 ;
     RECT 4.37000000 2.47700000 4.59000000 2.69700000 ;
     RECT 5.49000000 2.47700000 5.71000000 2.69700000 ;
     RECT 1.01000000 2.88200000 1.23000000 3.10200000 ;
     RECT 2.13000000 2.88200000 2.35000000 3.10200000 ;
     RECT 3.25000000 2.88200000 3.47000000 3.10200000 ;
     RECT 4.37000000 2.88200000 4.59000000 3.10200000 ;
     RECT 5.49000000 2.88200000 5.71000000 3.10200000 ;

    LAYER pdiffc ;
     RECT 0.45000000 3.28700000 0.67000000 3.50700000 ;
     RECT 6.05000000 3.55700000 6.27000000 3.77700000 ;
     RECT 1.57000000 4.50200000 1.79000000 4.72200000 ;

    LAYER ndiffc ;
     RECT 0.45000000 0.31700000 0.67000000 0.53700000 ;
     RECT 2.69000000 0.58700000 2.91000000 0.80700000 ;
     RECT 4.93000000 0.58700000 5.15000000 0.80700000 ;
     RECT 1.57000000 1.26200000 1.79000000 1.48200000 ;
     RECT 3.81000000 1.26200000 4.03000000 1.48200000 ;
     RECT 6.05000000 1.26200000 6.27000000 1.48200000 ;
     RECT 2.69000000 1.93700000 2.91000000 2.15700000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 6.72000000 0.24000000 ;
     RECT 0.37000000 0.24000000 0.75000000 0.61700000 ;
     RECT 2.61000000 0.50700000 2.99000000 0.88700000 ;
     RECT 4.85000000 0.50700000 5.23000000 0.88700000 ;
     RECT 1.49000000 1.18200000 1.87000000 1.56200000 ;
     RECT 3.73000000 1.18200000 4.11000000 1.56200000 ;
     RECT 5.97000000 1.18200000 6.35000000 1.56200000 ;
     RECT 2.61000000 1.85700000 2.99000000 2.23700000 ;
     RECT 5.41000000 2.39700000 5.79000000 2.77700000 ;
     RECT 0.93000000 2.39700000 1.31000000 2.47200000 ;
     RECT 1.49000000 2.39700000 1.87000000 2.47200000 ;
     RECT 0.93000000 2.47200000 1.87000000 2.70200000 ;
     RECT 1.49000000 2.70200000 1.87000000 2.77700000 ;
     RECT 0.93000000 2.70200000 1.31000000 3.18200000 ;
     RECT 3.73000000 2.12700000 4.11000000 2.20200000 ;
     RECT 3.24500000 2.20200000 4.11000000 2.39700000 ;
     RECT 3.17000000 2.39700000 4.11000000 2.43200000 ;
     RECT 3.73000000 2.43200000 4.11000000 2.50700000 ;
     RECT 3.17000000 2.43200000 3.55000000 3.18200000 ;
     RECT 4.29000000 2.39700000 4.67000000 3.18200000 ;
     RECT 5.41000000 2.80200000 5.79000000 3.18200000 ;
     RECT 1.49000000 3.07200000 1.87000000 3.14700000 ;
     RECT 2.05000000 2.39700000 2.43000000 3.14700000 ;
     RECT 1.49000000 3.14700000 2.43000000 3.18200000 ;
     RECT 1.49000000 3.18200000 2.35500000 3.37700000 ;
     RECT 1.49000000 3.37700000 1.87000000 3.45200000 ;
     RECT 0.37000000 3.20700000 0.75000000 3.58700000 ;
     RECT 5.97000000 3.47700000 6.35000000 3.85700000 ;
     RECT 1.49000000 4.42200000 1.87000000 4.80000000 ;
     RECT 0.00000000 4.80000000 6.72000000 5.28000000 ;

    LAYER via1 ;
     RECT 2.67000000 0.56700000 2.93000000 0.82700000 ;
     RECT 4.91000000 0.56700000 5.17000000 0.82700000 ;
     RECT 1.55000000 1.24200000 1.81000000 1.50200000 ;
     RECT 3.79000000 1.24200000 4.05000000 1.50200000 ;
     RECT 6.03000000 1.24200000 6.29000000 1.50200000 ;
     RECT 2.67000000 1.91700000 2.93000000 2.17700000 ;
     RECT 3.79000000 2.18700000 4.05000000 2.44700000 ;
     RECT 1.55000000 2.45700000 1.81000000 2.71700000 ;
     RECT 5.47000000 2.45700000 5.73000000 2.71700000 ;
     RECT 4.35000000 2.86200000 4.61000000 3.12200000 ;
     RECT 5.47000000 2.86200000 5.73000000 3.12200000 ;
     RECT 1.55000000 3.13200000 1.81000000 3.39200000 ;
     RECT 0.43000000 3.26700000 0.69000000 3.52700000 ;
     RECT 6.03000000 3.53700000 6.29000000 3.79700000 ;

    LAYER met2 ;
     RECT 2.61000000 0.50700000 2.99000000 0.55700000 ;
     RECT 4.85000000 0.50700000 5.23000000 0.55700000 ;
     RECT 2.61000000 0.55700000 5.23000000 0.83700000 ;
     RECT 2.61000000 0.83700000 2.99000000 0.88700000 ;
     RECT 4.85000000 0.83700000 5.23000000 0.88700000 ;
     RECT 3.73000000 2.12700000 4.11000000 2.50700000 ;
     RECT 1.49000000 2.39700000 1.87000000 2.77700000 ;
     RECT 4.29000000 2.80200000 4.67000000 3.18200000 ;
     RECT 5.41000000 2.39700000 5.79000000 3.18200000 ;
     RECT 1.49000000 3.07200000 1.87000000 3.45200000 ;
     RECT 1.49000000 1.18200000 1.87000000 1.23200000 ;
     RECT 3.73000000 1.18200000 4.11000000 1.23200000 ;
     RECT 5.97000000 1.18200000 6.35000000 1.23200000 ;
     RECT 0.42000000 1.23200000 6.35000000 1.51200000 ;
     RECT 1.49000000 1.51200000 1.87000000 1.56200000 ;
     RECT 3.73000000 1.51200000 4.11000000 1.56200000 ;
     RECT 5.97000000 1.51200000 6.35000000 1.56200000 ;
     RECT 0.42000000 1.51200000 0.70000000 3.20700000 ;
     RECT 0.37000000 3.20700000 0.75000000 3.58700000 ;
     RECT 2.61000000 1.85700000 2.99000000 2.23700000 ;
     RECT 2.66000000 2.23700000 2.94000000 3.52700000 ;
     RECT 5.97000000 3.47700000 6.35000000 3.52700000 ;
     RECT 2.66000000 3.52700000 6.35000000 3.80700000 ;
     RECT 5.97000000 3.80700000 6.35000000 3.85700000 ;

 END
END OAI41
