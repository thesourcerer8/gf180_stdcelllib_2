VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO AAAAOI3332
  CLASS CORE ;
  FOREIGN AAAAOI3332 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.550 BY 5.050 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.800 14.550 5.300 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.250 14.550 0.250 ;
    END
  END VGND
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 0.350 4.350 0.750 4.400 ;
        RECT 2.600 4.350 3.000 4.400 ;
        RECT 0.350 4.050 3.000 4.350 ;
        RECT 0.350 4.000 0.750 4.050 ;
        RECT 2.600 4.000 3.000 4.050 ;
    END
  END Y
  PIN C2
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 11.000 2.400 11.400 2.800 ;
    END
  END C2
  PIN A1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 2.050 2.400 2.450 2.800 ;
    END
  END A1
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 0.950 2.400 1.300 2.800 ;
    END
  END A
  PIN A2
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 3.150 2.400 3.550 2.800 ;
    END
  END A2
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 6.550 2.400 6.900 2.800 ;
    END
  END B
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 12.700 1.850 13.050 2.250 ;
        RECT 7.650 1.500 8.050 1.550 ;
        RECT 12.750 1.500 13.000 1.850 ;
        RECT 7.650 1.250 13.000 1.500 ;
        RECT 7.650 1.200 8.050 1.250 ;
    END
  END C
  PIN B2
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 4.300 2.400 4.650 2.800 ;
    END
  END B2
  PIN B1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 5.400 2.400 5.800 2.800 ;
    END
  END B1
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 9.900 2.400 10.250 2.800 ;
    END
  END D1
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 8.750 2.550 9.150 2.900 ;
    END
  END D
  PIN C1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 12.150 2.550 12.500 2.900 ;
    END
  END C1
END AAAAOI3332
END LIBRARY

