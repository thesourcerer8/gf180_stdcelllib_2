VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OAI41
  CLASS CORE ;
  FOREIGN OAI41 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.700 BY 5.050 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.800 6.700 5.300 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.250 6.700 0.250 ;
    END
  END VGND
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 2.600 0.850 3.000 0.900 ;
        RECT 4.850 0.850 5.250 0.900 ;
        RECT 2.600 0.550 5.250 0.850 ;
        RECT 2.600 0.500 3.000 0.550 ;
        RECT 4.850 0.500 5.250 0.550 ;
    END
  END Y
  PIN A1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 4.300 2.800 4.650 3.200 ;
    END
  END A1
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 1.500 2.400 1.850 2.800 ;
    END
  END B
  PIN A3
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 1.500 3.050 1.850 3.450 ;
    END
  END A3
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 5.400 2.400 5.800 3.200 ;
    END
  END A
  PIN A2
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 3.750 2.150 4.100 2.500 ;
    END
  END A2
END OAI41
END LIBRARY

